module  msrv32_pc_mux(input rst_in,
input [1:0] pc_src_in,
input [31:0] epc_in,
input [31:0] trap_address_in,
input branch_taken_in,
input [31:1] iaddr_in,
input ahb_ready_in,
input [31:0] pc_in,
output [31:0] iaddr_out,
output [31:0] pc_plus_4_out,
output misaligned_instr_out,
output reg [31:0] pc_mux_out);
reg [31:0] i_addr;
parameter BOOT_ADDRESS = 0;
wire [31:0] next_pc;
wire [31:0] w;
assign misaligned_instr_out=branch_taken_in & next_pc[1];
assign pc_plus_4_out=pc_in+32'h00000004;
assign next_pc=branch_taken_in?{iaddr_in,1'b0}:pc_plus_4_out;
assign w=ahb_ready_in?pc_mux_out:iaddr_out;
assign iaddr_out=rst_in?BOOT_ADDRESS:w;

always @(*)
 begin
case (pc_src_in)
2'b00:pc_mux_out=BOOT_ADDRESS;
2'b01:pc_mux_out=epc_in;
2'b10:pc_mux_out=trap_address_in;
2'b11:pc_mux_out=next_pc;
default : pc_mux_out = next_pc;

endcase
end

endmodule

